// q_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module q_sys (
    input  wire        clk_50_clk,                 //     clk_50.clk
    input  wire        clk_smc_clk,                //    clk_smc.clk
    output wire [13:0] memory_smc_mem_a,           // memory_smc.mem_a
    output wire [2:0]  memory_smc_mem_ba,          //           .mem_ba
    output wire [0:0]  memory_smc_mem_ck,          //           .mem_ck
    output wire [0:0]  memory_smc_mem_ck_n,        //           .mem_ck_n
    output wire [0:0]  memory_smc_mem_cke,         //           .mem_cke
    output wire [0:0]  memory_smc_mem_cs_n,        //           .mem_cs_n
    output wire [7:0]  memory_smc_mem_dm,          //           .mem_dm
    output wire [0:0]  memory_smc_mem_ras_n,       //           .mem_ras_n
    output wire [0:0]  memory_smc_mem_cas_n,       //           .mem_cas_n
    output wire [0:0]  memory_smc_mem_we_n,        //           .mem_we_n
    output wire        memory_smc_mem_reset_n,     //           .mem_reset_n
    inout  wire [63:0] memory_smc_mem_dq,          //           .mem_dq
    inout  wire [7:0]  memory_smc_mem_dqs,         //           .mem_dqs
    inout  wire [7:0]  memory_smc_mem_dqs_n,       //           .mem_dqs_n
    output wire [0:0]  memory_smc_mem_odt,         //           .mem_odt
    input  wire        oct_hmc_rzqin,              //    oct_hmc.rzqin
    input  wire        reset_50_reset_n,           //   reset_50.reset_n
    input  wire        reset_smc_reset_n,          //  reset_smc.reset_n
    output wire        smc_error_mon,              //        smc.error_mon
    output wire        smc_status_mon,             //           .status_mon
    output wire        smc_status_cal_fail_mon,    // smc_status.cal_fail_mon
    output wire        smc_status_cal_success_mon, //           .cal_success_mon
    output wire        smc_status_init_done_mon,   //           .init_done_mon
    input  wire        tg_smc_reset_n,              //     tg_smc.reset_n
    
    output wire         avl_ready,        
    input  wire         avl_burstbegin,       
    input  wire [24:0]  avl_addr,             
    output wire         avl_rdata_valid,      
    output wire [255:0] avl_rdata,            
    input  wire [255:0] avl_wdata,        
    input  wire         avl_read_req,     
    input  wire         avl_write_req,    
    input  wire [9:0]   avl_size,         
    output wire         local_init_done,  
    output wire         local_cal_success,
    output wire         local_cal_fail,
    
    output wire         afi_clk
    
);

	wire  [15:0] hmc_0_fpga_sdram_oct_sharing_parallelterminationcontrol;    // hmc_0:fpga_sdram_oct_sharing_parallelterminationcontrol
	wire  [15:0] hmc_0_fpga_sdram_oct_sharing_seriesterminationcontrol;      // hmc_0:fpga_sdram_oct_sharing_seriesterminationcontrol
    
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out

                      
    
	altera_mem_if_oct_cyclonev #(
		.OCT_TERM_CONTROL_WIDTH (16)
	) oct0 (
		.oct_rzqin                  (oct_hmc_rzqin),                                           //         oct.rzqin
		.seriesterminationcontrol   (hmc_0_fpga_sdram_oct_sharing_seriesterminationcontrol),   // oct_sharing.seriesterminationcontrol
		.parallelterminationcontrol (hmc_0_fpga_sdram_oct_sharing_parallelterminationcontrol)  //            .parallelterminationcontrol
        );

	q_sys_smc_0 smc_0 (
		.memory_mem_a                                              (memory_smc_mem_a),           //                             memory.mem_a
		.memory_mem_ba                                             (memory_smc_mem_ba),          //                                   .mem_ba
		.memory_mem_ck                                             (memory_smc_mem_ck),          //                                   .mem_ck
		.memory_mem_ck_n                                           (memory_smc_mem_ck_n),        //                                   .mem_ck_n
		.memory_mem_cke                                            (memory_smc_mem_cke),         //                                   .mem_cke
		.memory_mem_cs_n                                           (memory_smc_mem_cs_n),        //                                   .mem_cs_n
		.memory_mem_dm                                             (memory_smc_mem_dm),          //                                   .mem_dm
		.memory_mem_ras_n                                          (memory_smc_mem_ras_n),       //                                   .mem_ras_n
		.memory_mem_cas_n                                          (memory_smc_mem_cas_n),       //                                   .mem_cas_n
		.memory_mem_we_n                                           (memory_smc_mem_we_n),        //                                   .mem_we_n
		.memory_mem_reset_n                                        (memory_smc_mem_reset_n),     //                                   .mem_reset_n
		.memory_mem_dq                                             (memory_smc_mem_dq),          //                                   .mem_dq
		.memory_mem_dqs                                            (memory_smc_mem_dqs),         //                                   .mem_dqs
		.memory_mem_dqs_n                                          (memory_smc_mem_dqs_n),       //                                   .mem_dqs_n
		.memory_mem_odt                                            (memory_smc_mem_odt),         //                                   .mem_odt
		.clk_100_clk                                               (clk_smc_clk),                //                            clk_100.clk
		.clk_50_clk                                                (clk_50_clk),                 //                             clk_50.clk
		.reset_50_reset_n                                          (reset_50_reset_n),           //                           reset_50.reset_n
		.master_driver_msgdma_0_conduit_end_error_mon              (smc_error_mon),              // master_driver_msgdma_0_conduit_end.error_mon
		.master_driver_msgdma_0_conduit_end_status_mon             (smc_status_mon),             //                                   .status_mon
		.msgdma_0_status_mon_out_cal_fail_mon                      (smc_status_cal_fail_mon),    //            msgdma_0_status_mon_out.cal_fail_mon
		.msgdma_0_status_mon_out_cal_success_mon                   (smc_status_cal_success_mon), //                                   .cal_success_mon
		.msgdma_0_status_mon_out_init_done_mon                     (smc_status_init_done_mon),   //                                   .init_done_mon
        
        .avl_ready          (avl_ready),        
        .avl_burstbegin     (avl_burstbegin),   
        .avl_addr           (avl_addr),         
        .avl_rdata_valid    (avl_rdata_valid),  
        .avl_rdata          (avl_rdata),        
        .avl_wdata          (avl_wdata),        
        .avl_read_req       (avl_read_req),     
        .avl_write_req      (avl_write_req),    
        .avl_size           (avl_size),         
        .local_init_done    (local_init_done),  
        .local_cal_success  (local_cal_success),
        .local_cal_fail     (local_cal_fail),   
		  
		 .afi_clk            (afi_clk),
        
		.mem_if_ddr3_emif_0_oct_sharing_seriesterminationcontrol   (hmc_0_fpga_sdram_oct_sharing_seriesterminationcontrol),   //     mem_if_ddr3_emif_0_oct_sharing.seriesterminationcontrol
		.mem_if_ddr3_emif_0_oct_sharing_parallelterminationcontrol (hmc_0_fpga_sdram_oct_sharing_parallelterminationcontrol), //                                   .parallelterminationcontrol
		.tg_reset_n                                                (tg_smc_reset_n),                                          //                                 tg.reset_n
		.reset_reset_n                                             (reset_smc_reset_n)                                        //                              reset.reset_n
	);

	/*altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_50_reset_n),              // reset_in0.reset
		.clk            (clk_50_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset) // reset_out.reset
		.reset_req      ().                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);*/

endmodule
