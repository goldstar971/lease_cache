//`include "riscv.h"

module stage1_instruction_decode(

	input 	[31:0]	instruction_i,
	output 	[15:0]	encoding_o, 		// one hot encoding of instruction type
	output 	[6:0] 	func7_o,
	output 	[2:0] 	func3_o,
	output   [4:0] fsrc3_o,
	output 	[4:0]	fsrc2_o,
	output 	[4:0]	fsrc1_o,
	output 	[4:0]	fdest_o,
	output   [4:0] func5_o,
	output   [2:0] rm_o,
	output 	[31:0]	imm32_o, 			// generate immediate value during decode because 32b imm is consistent across all 32b extensions
	output 			exception_o 		// unknown opcode

);

// port mappings
// -----------------------------------------------------------------------------------
reg 	[15:0]	encoding_reg;
reg 	[6:0] 	func7_reg;
reg 	[2:0] 	func3_reg;
reg   [4:0]   func5_reg;
reg   [2:0]   rm_reg;
reg 	[4:0]	fsrc2_reg;
reg 	[4:0]	fsrc3_reg;
reg 	[4:0]	fsrc1_reg;
reg 	[4:0]	fdest_reg;
reg 	[31:0]	imm32_reg;
reg 			exception_reg;

assign encoding_o 	= encoding_reg;
assign func7_o 		= func7_reg;
assign func5_o 		= func5_reg;
assign func3_o 		= func3_reg;
assign fsrc2_o 		= fsrc2_reg;
assign fsrc1_o 		= fsrc1_reg;
assign fdest_o 		= fdest_reg;
assign imm32_o 		= imm32_reg;
assign fsrc3_o 		= fsrc3_reg;
assign rm_o  			=	  rm_reg;
assign exception_o 	= exception_reg;


// stage combinational logic
// -----------------------------------------------------------------------------------

always @(*) begin

	// default outputs
	// -------------------------------------------------------------------------------
	encoding_reg 	= `ENCODING_NONE;
	func7_reg  		= 'b0;
	func5_reg      = 'b0;
	func3_reg  		= 'b0;
	fsrc3_reg      = 'b0;
	fsrc2_reg  		= 'b0;
	fsrc1_reg  		= 'b0;
	fdest_reg  		= 'b0;
	imm32_reg  		= 'b0;
	rm_reg 			= 'b0;
	exception_reg 	= 1'b0;

	// instruction decoding - by opcode field
	// -------------------------------------------------------------------------------
	case(instruction_i[6:0])

		// RV32I extension instructions
		// ---------------------------------------------------------------------------
		// supported instructions
		`RV32I_OPCODE_LUI: begin
			encoding_reg 	= `ENCODING_LUI;		
			fdest_reg 		= instruction_i[11:7];
			imm32_reg 		= {instruction_i[31:12],12'h000};
		end

		`RV32I_OPCODE_AUIPC: begin
			encoding_reg 	= `ENCODING_AUIPC;		
			fdest_reg 		= instruction_i[11:7];
			imm32_reg 		= {instruction_i[31:12],12'h000};
		end

		`RV32I_OPCODE_JAL: 	begin												
			encoding_reg 	= `ENCODING_JAL;		
			fdest_reg 		= instruction_i[11:7];
			imm32_reg 		= {{11{instruction_i[31]}}, instruction_i[31], instruction_i[19:12], instruction_i[20], instruction_i[30:21], 1'b0};
		end

		`RV32I_OPCODE_JALR: begin
			encoding_reg 	= `ENCODING_JALR;
			fsrc1_reg 		= instruction_i[19:15];
			fdest_reg 		= instruction_i[11:7];
			imm32_reg 		= {{20{instruction_i[31]}},instruction_i[31:20]};
		end

		`RV32I_OPCODE_LOAD: begin
			encoding_reg 	= `ENCODING_LOAD;
			fsrc1_reg 		= instruction_i[19:15];
			func3_reg 		= instruction_i[14:12];
			fdest_reg 		= instruction_i[11:7];
			imm32_reg 		= {{20{instruction_i[31]}},instruction_i[31:20]};
		end 

		`RV32I_OPCODE_ARITH_IMM: begin
			encoding_reg 	= `ENCODING_ARITH_IMM;
			fsrc1_reg 		= instruction_i[19:15];
			func3_reg 		= instruction_i[14:12];
			fdest_reg 		= instruction_i[11:7];
			imm32_reg 		= {{20{instruction_i[31]}},instruction_i[31:20]};
		end

		`RV32I_OPCODE_BRANCH: begin
			encoding_reg 	= `ENCODING_BRANCH;
			fsrc2_reg 		= instruction_i[24:20]; 
			fsrc1_reg 		= instruction_i[19:15]; 
			func3_reg 		= instruction_i[14:12];
			imm32_reg 		= {{19{instruction_i[31]}},instruction_i[31],instruction_i[7],instruction_i[30:25],instruction_i[11:8],1'b0};
		end

		`RV32I_OPCODE_STORE: begin
			encoding_reg 	= `ENCODING_STORE;
			fsrc2_reg 		= instruction_i[24:20]; 
			fsrc1_reg 		= instruction_i[19:15]; 
			func3_reg 		= instruction_i[14:12];
			imm32_reg 		= {{20{instruction_i[31]}},instruction_i[31:25],instruction_i[11:7]};
		end
		


		// RV32I register-register and RV32M extension instructions
		// ---------------------------------------------------------------------------
		`RV32I_OPCODE_ARITH_REG: begin
			encoding_reg = `ENCODING_ARITH_REG;
			{func7_reg,fsrc2_reg,fsrc1_reg,func3_reg,fdest_reg} = instruction_i[31:7];
		end
		
		
		//RV32F single precision extension instructions
		`RV32F_OPCODE_LOAD: begin
			encoding_reg =`ENCODING_FLOAD;
			{fsrc1_reg,fdest_reg,imm32_reg}={instruction_i[19:15],instruction_i[11:7],
			{20{instruction_i[31]}},instruction_i[31:20]}; 
		end
		`RV32F_OPCODE_STORE: begin
			encoding_reg=`ENCODING_FSTORE;
			{fsrc2_reg,fsrc1_reg,imm32_reg}={instruction_i[24:20],instruction_i[19:15],
			{{20{instruction_i[31]}},instruction_i[31:25],instruction_i[11:7]}}; 
		end
		`RV32F_OPCODE_FMADD: begin
			encoding_reg =`ENCODING_FMADD;
			{fsrc1_reg,fsrc2_reg,fdest_reg,rm_reg,fsrc3_reg}={instruction_i[19:15],
			instruction_i[24:20],instruction_i[11:7],instruction_i[14:12],instruction_i[31:27]};
		end
			`RV32F_OPCODE_FMSUB: begin
			encoding_reg =`ENCODING_FMSUB;
			{fsrc1_reg,fsrc2_reg,fdest_reg,rm_reg,fsrc3_reg}={instruction_i[19:15],
			instruction_i[24:20],instruction_i[11:7],instruction_i[14:12],instruction_i[31:27]};
		end
			`RV32F_OPCODE_FNMADD: begin
			encoding_reg =`ENCODING_FNMADD;
			{fsrc1_reg,fsrc2_reg,fdest_reg,rm_reg,fsrc3_reg}={instruction_i[19:15]
			,instruction_i[24:20],instruction_i[11:7],instruction_i[14:12],instruction_i[31:27]};
		end
			`RV32F_OPCODE_FNMSUB: begin
			encoding_reg =`ENCODING_FNMSUB;
			{fsrc1_reg,fsrc2_reg,fdest_reg,rm_reg,fsrc3_reg}={instruction_i[19:15]
			,instruction_i[24:20],instruction_i[11:7],instruction_i[14:12],instruction_i[31:27]};
		end
		`RV32F_OPCODE_ARITH: begin
			encoding_reg =`ENCODING_FARITH;
			{fsrc1_reg,fsrc2_reg,fdest_reg,rm_reg,func5_reg}={instruction_i[19:15]
			,instruction_i[24:20],instruction_i[11:7],instruction_i[14:12],instruction_i[31:27]};
		end
		// Unknown instructions - raise exception
		// ---------------------------------------------------------------------------
		default: begin
			exception_reg 	= 1'b1;
		end

	endcase

end

endmodule