// q_sys_smc_0.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module q_sys_smc_0 (
		output wire [13:0] memory_mem_a,         
		output wire [2:0]  memory_mem_ba,        
		output wire [0:0]  memory_mem_ck,        
		output wire [0:0]  memory_mem_ck_n,      
		output wire [0:0]  memory_mem_cke,       
		output wire [0:0]  memory_mem_cs_n,      
		output wire [7:0]  memory_mem_dm,        
		output wire [0:0]  memory_mem_ras_n,     
		output wire [0:0]  memory_mem_cas_n,     
		output wire [0:0]  memory_mem_we_n,      
		output wire        memory_mem_reset_n,   
		inout  wire [63:0] memory_mem_dq,        
		inout  wire [7:0]  memory_mem_dqs,       
		inout  wire [7:0]  memory_mem_dqs_n,     
		output wire [0:0]  memory_mem_odt,       
        
        output wire         avl_ready,        
        input  wire         avl_burstbegin,   
        input  wire [24:0]  avl_addr,         
        output wire         avl_rdata_valid,  
        output wire [255:0] avl_rdata,        
        input  wire [255:0] avl_wdata,        
        input  wire         avl_read_req,     
        input  wire         avl_write_req,    
        input  wire [9:0]   avl_size,         
        output wire         local_init_done,  
        output wire         local_cal_success,
        output wire         local_cal_fail,   
		
		  output wire 	       afi_clk,
          
        /*output wire risc_50_clk,
        output wire risc_40_clk,
        output wire risc_30_clk,
        output wire risc_20_clk,
        output wire risc_10_clk,*/
        
		input  wire        clk_100,     
		//input 	clk_phy_100,                                        //                            clk_100.clk

		input  wire [15:0] seriesterminationcontrol,   //     mem_if_ddr3_emif_0_oct_sharing.seriesterminationcontrol
		input  wire [15:0] parallelterminationcontrol, //                                   .parallelterminationcontrol
		input  wire        reset_n                                              //                              reset.reset_n
	);

	q_sys_smc_0_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk                (clk_100),                    //      pll_ref_clk.clk
		.global_reset_n             (reset_n),                  //     global_reset.reset_n
		.soft_reset_n               (reset_n),                  //       soft_reset.reset_n
		.afi_clk                    (afi_clk), //          afi_clk.clk
		.afi_half_clk               (),                               //     afi_half_clk.clk
		.afi_reset_n                (),                               //        afi_reset.reset_n
		.afi_reset_export_n         (),                               // afi_reset_export.reset_n
		.mem_a                      (memory_mem_a),                   //           memory.mem_a
		.mem_ba                     (memory_mem_ba),                  //                 .mem_ba
		.mem_ck                     (memory_mem_ck),                  //                 .mem_ck
		.mem_ck_n                   (memory_mem_ck_n),                //                 .mem_ck_n
		.mem_cke                    (memory_mem_cke),                 //                 .mem_cke
		.mem_cs_n                   (memory_mem_cs_n),                //                 .mem_cs_n
		.mem_dm                     (memory_mem_dm),                  //                 .mem_dm
		.mem_ras_n                  (memory_mem_ras_n),               //                 .mem_ras_n
		.mem_cas_n                  (memory_mem_cas_n),               //                 .mem_cas_n
		.mem_we_n                   (memory_mem_we_n),                //                 .mem_we_n
		.mem_reset_n                (memory_mem_reset_n),             //                 .mem_reset_n
		.mem_dq                     (memory_mem_dq),                  //                 .mem_dq
		.mem_dqs                    (memory_mem_dqs),                 //                 .mem_dqs
		.mem_dqs_n                  (memory_mem_dqs_n),               //                 .mem_dqs_n
		.mem_odt                    (memory_mem_odt),                 //                 .mem_odt
		.avl_ready                  (avl_ready),             //     avl.waitrequest_n
		.avl_burstbegin             (avl_burstbegin),        //    .beginbursttransfer
		.avl_addr                   (avl_addr),              //    .address
		.avl_rdata_valid            (avl_rdata_valid),       //    .readdatavalid
		.avl_rdata                  (avl_rdata),             //    .readdata
		.avl_wdata                  (avl_wdata),             //    .writedata
		.avl_read_req               (avl_read_req),          //    .read
		.avl_write_req              (avl_write_req),         //    .write
		.avl_size                   (avl_size),              //    .burstcount
		.local_init_done            (local_init_done),       //     status.local_init_done
		.local_cal_success          (local_cal_success),     //    .local_cal_success
		.local_cal_fail             (local_cal_fail),        //    .local_cal_fail
		.seriesterminationcontrol   (seriesterminationcontrol),     //      oct_sharing.seriesterminationcontrol
		.parallelterminationcontrol (parallelterminationcontrol),   //                 .parallelterminationcontrol
		.pll_mem_clk                (),                                                            //      pll_sharing.pll_mem_clk
		.pll_write_clk              (),                                                            //                 .pll_write_clk
		.pll_locked                 (),                                                            //                 .pll_locked
		.pll_write_clk_pre_phy_clk  (),                                                            //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (),                                                            //                 .pll_addr_cmd_clk
		.pll_avl_clk                (),                                                            //                 .pll_avl_clk
		.pll_config_clk             (),                                                            //                 .pll_config_clk
		.pll_mem_phy_clk            (),                                                            //                 .pll_mem_phy_clk
		.afi_phy_clk                (),                                                            //                 .afi_phy_clk
		.pll_avl_phy_clk            ()                                                             //                 .pll_avl_phy_clk
        
        /*.risc_50_clk                (risc_50_clk),
        .risc_40_clk                (risc_40_clk),
        .risc_30_clk                (risc_30_clk),
        .risc_20_clk                (risc_20_clk),
        .risc_10_clk                (risc_10_clk)*/
	);



endmodule
