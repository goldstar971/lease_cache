module eviction_bit_tracker #(
	parameter N_LINES 	= 0,
	parameter BINS 		= 0
)(
	input 
);

// parameterizations
// ---------------------------------------------------
localparam BW_LINES = `CLOG2(N_LINES);



endmodule