module tag_match_encoder_9b(
input [511:0] match_bits,
	output reg [8:0] match_index_reg,
 output reg actual_match);
wire [31:0] or_o[8:0];
wire [8:0] match_index;
	assign or_o[0][0]=|({match_bits[1],match_bits[3],match_bits[5],match_bits[7],match_bits[9],match_bits[11],match_bits[13],match_bits[15]});
	assign or_o[0][1]=|({match_bits[17],match_bits[19],match_bits[21],match_bits[23],match_bits[25],match_bits[27],match_bits[29],match_bits[31]});
	assign or_o[0][2]=|({match_bits[33],match_bits[35],match_bits[37],match_bits[39],match_bits[41],match_bits[43],match_bits[45],match_bits[47]});
	assign or_o[0][3]=|({match_bits[49],match_bits[51],match_bits[53],match_bits[55],match_bits[57],match_bits[59],match_bits[61],match_bits[63]});
	assign or_o[0][4]=|({match_bits[65],match_bits[67],match_bits[69],match_bits[71],match_bits[73],match_bits[75],match_bits[77],match_bits[79]});
	assign or_o[0][5]=|({match_bits[81],match_bits[83],match_bits[85],match_bits[87],match_bits[89],match_bits[91],match_bits[93],match_bits[95]});
	assign or_o[0][6]=|({match_bits[97],match_bits[99],match_bits[101],match_bits[103],match_bits[105],match_bits[107],match_bits[109],match_bits[111]});
	assign or_o[0][7]=|({match_bits[113],match_bits[115],match_bits[117],match_bits[119],match_bits[121],match_bits[123],match_bits[125],match_bits[127]});
	assign or_o[0][8]=|({match_bits[129],match_bits[131],match_bits[133],match_bits[135],match_bits[137],match_bits[139],match_bits[141],match_bits[143]});
	assign or_o[0][9]=|({match_bits[145],match_bits[147],match_bits[149],match_bits[151],match_bits[153],match_bits[155],match_bits[157],match_bits[159]});
	assign or_o[0][10]=|({match_bits[161],match_bits[163],match_bits[165],match_bits[167],match_bits[169],match_bits[171],match_bits[173],match_bits[175]});
	assign or_o[0][11]=|({match_bits[177],match_bits[179],match_bits[181],match_bits[183],match_bits[185],match_bits[187],match_bits[189],match_bits[191]});
	assign or_o[0][12]=|({match_bits[193],match_bits[195],match_bits[197],match_bits[199],match_bits[201],match_bits[203],match_bits[205],match_bits[207]});
	assign or_o[0][13]=|({match_bits[209],match_bits[211],match_bits[213],match_bits[215],match_bits[217],match_bits[219],match_bits[221],match_bits[223]});
	assign or_o[0][14]=|({match_bits[225],match_bits[227],match_bits[229],match_bits[231],match_bits[233],match_bits[235],match_bits[237],match_bits[239]});
	assign or_o[0][15]=|({match_bits[241],match_bits[243],match_bits[245],match_bits[247],match_bits[249],match_bits[251],match_bits[253],match_bits[255]});
	assign or_o[0][16]=|({match_bits[257],match_bits[259],match_bits[261],match_bits[263],match_bits[265],match_bits[267],match_bits[269],match_bits[271]});
	assign or_o[0][17]=|({match_bits[273],match_bits[275],match_bits[277],match_bits[279],match_bits[281],match_bits[283],match_bits[285],match_bits[287]});
	assign or_o[0][18]=|({match_bits[289],match_bits[291],match_bits[293],match_bits[295],match_bits[297],match_bits[299],match_bits[301],match_bits[303]});
	assign or_o[0][19]=|({match_bits[305],match_bits[307],match_bits[309],match_bits[311],match_bits[313],match_bits[315],match_bits[317],match_bits[319]});
	assign or_o[0][20]=|({match_bits[321],match_bits[323],match_bits[325],match_bits[327],match_bits[329],match_bits[331],match_bits[333],match_bits[335]});
	assign or_o[0][21]=|({match_bits[337],match_bits[339],match_bits[341],match_bits[343],match_bits[345],match_bits[347],match_bits[349],match_bits[351]});
	assign or_o[0][22]=|({match_bits[353],match_bits[355],match_bits[357],match_bits[359],match_bits[361],match_bits[363],match_bits[365],match_bits[367]});
	assign or_o[0][23]=|({match_bits[369],match_bits[371],match_bits[373],match_bits[375],match_bits[377],match_bits[379],match_bits[381],match_bits[383]});
	assign or_o[0][24]=|({match_bits[385],match_bits[387],match_bits[389],match_bits[391],match_bits[393],match_bits[395],match_bits[397],match_bits[399]});
	assign or_o[0][25]=|({match_bits[401],match_bits[403],match_bits[405],match_bits[407],match_bits[409],match_bits[411],match_bits[413],match_bits[415]});
	assign or_o[0][26]=|({match_bits[417],match_bits[419],match_bits[421],match_bits[423],match_bits[425],match_bits[427],match_bits[429],match_bits[431]});
	assign or_o[0][27]=|({match_bits[433],match_bits[435],match_bits[437],match_bits[439],match_bits[441],match_bits[443],match_bits[445],match_bits[447]});
	assign or_o[0][28]=|({match_bits[449],match_bits[451],match_bits[453],match_bits[455],match_bits[457],match_bits[459],match_bits[461],match_bits[463]});
	assign or_o[0][29]=|({match_bits[465],match_bits[467],match_bits[469],match_bits[471],match_bits[473],match_bits[475],match_bits[477],match_bits[479]});
	assign or_o[0][30]=|({match_bits[481],match_bits[483],match_bits[485],match_bits[487],match_bits[489],match_bits[491],match_bits[493],match_bits[495]});
	assign or_o[0][31]=|({match_bits[497],match_bits[499],match_bits[501],match_bits[503],match_bits[505],match_bits[507],match_bits[509],match_bits[511]});
	assign match_index[0]=|({or_o[0][0],or_o[0][1],or_o[0][2],or_o[0][3],or_o[0][4],or_o[0][5],or_o[0][6],or_o[0][7],or_o[0][8],or_o[0][9],or_o[0][10],or_o[0][11],or_o[0][12],or_o[0][13],or_o[0][14],or_o[0][15],or_o[0][16],or_o[0][17],or_o[0][18],or_o[0][19],or_o[0][20],or_o[0][21],or_o[0][22],or_o[0][23],or_o[0][24],or_o[0][25],or_o[0][26],or_o[0][27],or_o[0][28],or_o[0][29],or_o[0][30],or_o[0][31]});
	assign or_o[1][0]=|({match_bits[2],match_bits[3],match_bits[6],match_bits[7],match_bits[10],match_bits[11],match_bits[14],match_bits[15]});
	assign or_o[1][1]=|({match_bits[18],match_bits[19],match_bits[22],match_bits[23],match_bits[26],match_bits[27],match_bits[30],match_bits[31]});
	assign or_o[1][2]=|({match_bits[34],match_bits[35],match_bits[38],match_bits[39],match_bits[42],match_bits[43],match_bits[46],match_bits[47]});
	assign or_o[1][3]=|({match_bits[50],match_bits[51],match_bits[54],match_bits[55],match_bits[58],match_bits[59],match_bits[62],match_bits[63]});
	assign or_o[1][4]=|({match_bits[66],match_bits[67],match_bits[70],match_bits[71],match_bits[74],match_bits[75],match_bits[78],match_bits[79]});
	assign or_o[1][5]=|({match_bits[82],match_bits[83],match_bits[86],match_bits[87],match_bits[90],match_bits[91],match_bits[94],match_bits[95]});
	assign or_o[1][6]=|({match_bits[98],match_bits[99],match_bits[102],match_bits[103],match_bits[106],match_bits[107],match_bits[110],match_bits[111]});
	assign or_o[1][7]=|({match_bits[114],match_bits[115],match_bits[118],match_bits[119],match_bits[122],match_bits[123],match_bits[126],match_bits[127]});
	assign or_o[1][8]=|({match_bits[130],match_bits[131],match_bits[134],match_bits[135],match_bits[138],match_bits[139],match_bits[142],match_bits[143]});
	assign or_o[1][9]=|({match_bits[146],match_bits[147],match_bits[150],match_bits[151],match_bits[154],match_bits[155],match_bits[158],match_bits[159]});
	assign or_o[1][10]=|({match_bits[162],match_bits[163],match_bits[166],match_bits[167],match_bits[170],match_bits[171],match_bits[174],match_bits[175]});
	assign or_o[1][11]=|({match_bits[178],match_bits[179],match_bits[182],match_bits[183],match_bits[186],match_bits[187],match_bits[190],match_bits[191]});
	assign or_o[1][12]=|({match_bits[194],match_bits[195],match_bits[198],match_bits[199],match_bits[202],match_bits[203],match_bits[206],match_bits[207]});
	assign or_o[1][13]=|({match_bits[210],match_bits[211],match_bits[214],match_bits[215],match_bits[218],match_bits[219],match_bits[222],match_bits[223]});
	assign or_o[1][14]=|({match_bits[226],match_bits[227],match_bits[230],match_bits[231],match_bits[234],match_bits[235],match_bits[238],match_bits[239]});
	assign or_o[1][15]=|({match_bits[242],match_bits[243],match_bits[246],match_bits[247],match_bits[250],match_bits[251],match_bits[254],match_bits[255]});
	assign or_o[1][16]=|({match_bits[258],match_bits[259],match_bits[262],match_bits[263],match_bits[266],match_bits[267],match_bits[270],match_bits[271]});
	assign or_o[1][17]=|({match_bits[274],match_bits[275],match_bits[278],match_bits[279],match_bits[282],match_bits[283],match_bits[286],match_bits[287]});
	assign or_o[1][18]=|({match_bits[290],match_bits[291],match_bits[294],match_bits[295],match_bits[298],match_bits[299],match_bits[302],match_bits[303]});
	assign or_o[1][19]=|({match_bits[306],match_bits[307],match_bits[310],match_bits[311],match_bits[314],match_bits[315],match_bits[318],match_bits[319]});
	assign or_o[1][20]=|({match_bits[322],match_bits[323],match_bits[326],match_bits[327],match_bits[330],match_bits[331],match_bits[334],match_bits[335]});
	assign or_o[1][21]=|({match_bits[338],match_bits[339],match_bits[342],match_bits[343],match_bits[346],match_bits[347],match_bits[350],match_bits[351]});
	assign or_o[1][22]=|({match_bits[354],match_bits[355],match_bits[358],match_bits[359],match_bits[362],match_bits[363],match_bits[366],match_bits[367]});
	assign or_o[1][23]=|({match_bits[370],match_bits[371],match_bits[374],match_bits[375],match_bits[378],match_bits[379],match_bits[382],match_bits[383]});
	assign or_o[1][24]=|({match_bits[386],match_bits[387],match_bits[390],match_bits[391],match_bits[394],match_bits[395],match_bits[398],match_bits[399]});
	assign or_o[1][25]=|({match_bits[402],match_bits[403],match_bits[406],match_bits[407],match_bits[410],match_bits[411],match_bits[414],match_bits[415]});
	assign or_o[1][26]=|({match_bits[418],match_bits[419],match_bits[422],match_bits[423],match_bits[426],match_bits[427],match_bits[430],match_bits[431]});
	assign or_o[1][27]=|({match_bits[434],match_bits[435],match_bits[438],match_bits[439],match_bits[442],match_bits[443],match_bits[446],match_bits[447]});
	assign or_o[1][28]=|({match_bits[450],match_bits[451],match_bits[454],match_bits[455],match_bits[458],match_bits[459],match_bits[462],match_bits[463]});
	assign or_o[1][29]=|({match_bits[466],match_bits[467],match_bits[470],match_bits[471],match_bits[474],match_bits[475],match_bits[478],match_bits[479]});
	assign or_o[1][30]=|({match_bits[482],match_bits[483],match_bits[486],match_bits[487],match_bits[490],match_bits[491],match_bits[494],match_bits[495]});
	assign or_o[1][31]=|({match_bits[498],match_bits[499],match_bits[502],match_bits[503],match_bits[506],match_bits[507],match_bits[510],match_bits[511]});
	assign match_index[1]=|({or_o[1][0],or_o[1][1],or_o[1][2],or_o[1][3],or_o[1][4],or_o[1][5],or_o[1][6],or_o[1][7],or_o[1][8],or_o[1][9],or_o[1][10],or_o[1][11],or_o[1][12],or_o[1][13],or_o[1][14],or_o[1][15],or_o[1][16],or_o[1][17],or_o[1][18],or_o[1][19],or_o[1][20],or_o[1][21],or_o[1][22],or_o[1][23],or_o[1][24],or_o[1][25],or_o[1][26],or_o[1][27],or_o[1][28],or_o[1][29],or_o[1][30],or_o[1][31]});
	assign or_o[2][0]=|({match_bits[4],match_bits[5],match_bits[6],match_bits[7],match_bits[12],match_bits[13],match_bits[14],match_bits[15]});
	assign or_o[2][1]=|({match_bits[20],match_bits[21],match_bits[22],match_bits[23],match_bits[28],match_bits[29],match_bits[30],match_bits[31]});
	assign or_o[2][2]=|({match_bits[36],match_bits[37],match_bits[38],match_bits[39],match_bits[44],match_bits[45],match_bits[46],match_bits[47]});
	assign or_o[2][3]=|({match_bits[52],match_bits[53],match_bits[54],match_bits[55],match_bits[60],match_bits[61],match_bits[62],match_bits[63]});
	assign or_o[2][4]=|({match_bits[68],match_bits[69],match_bits[70],match_bits[71],match_bits[76],match_bits[77],match_bits[78],match_bits[79]});
	assign or_o[2][5]=|({match_bits[84],match_bits[85],match_bits[86],match_bits[87],match_bits[92],match_bits[93],match_bits[94],match_bits[95]});
	assign or_o[2][6]=|({match_bits[100],match_bits[101],match_bits[102],match_bits[103],match_bits[108],match_bits[109],match_bits[110],match_bits[111]});
	assign or_o[2][7]=|({match_bits[116],match_bits[117],match_bits[118],match_bits[119],match_bits[124],match_bits[125],match_bits[126],match_bits[127]});
	assign or_o[2][8]=|({match_bits[132],match_bits[133],match_bits[134],match_bits[135],match_bits[140],match_bits[141],match_bits[142],match_bits[143]});
	assign or_o[2][9]=|({match_bits[148],match_bits[149],match_bits[150],match_bits[151],match_bits[156],match_bits[157],match_bits[158],match_bits[159]});
	assign or_o[2][10]=|({match_bits[164],match_bits[165],match_bits[166],match_bits[167],match_bits[172],match_bits[173],match_bits[174],match_bits[175]});
	assign or_o[2][11]=|({match_bits[180],match_bits[181],match_bits[182],match_bits[183],match_bits[188],match_bits[189],match_bits[190],match_bits[191]});
	assign or_o[2][12]=|({match_bits[196],match_bits[197],match_bits[198],match_bits[199],match_bits[204],match_bits[205],match_bits[206],match_bits[207]});
	assign or_o[2][13]=|({match_bits[212],match_bits[213],match_bits[214],match_bits[215],match_bits[220],match_bits[221],match_bits[222],match_bits[223]});
	assign or_o[2][14]=|({match_bits[228],match_bits[229],match_bits[230],match_bits[231],match_bits[236],match_bits[237],match_bits[238],match_bits[239]});
	assign or_o[2][15]=|({match_bits[244],match_bits[245],match_bits[246],match_bits[247],match_bits[252],match_bits[253],match_bits[254],match_bits[255]});
	assign or_o[2][16]=|({match_bits[260],match_bits[261],match_bits[262],match_bits[263],match_bits[268],match_bits[269],match_bits[270],match_bits[271]});
	assign or_o[2][17]=|({match_bits[276],match_bits[277],match_bits[278],match_bits[279],match_bits[284],match_bits[285],match_bits[286],match_bits[287]});
	assign or_o[2][18]=|({match_bits[292],match_bits[293],match_bits[294],match_bits[295],match_bits[300],match_bits[301],match_bits[302],match_bits[303]});
	assign or_o[2][19]=|({match_bits[308],match_bits[309],match_bits[310],match_bits[311],match_bits[316],match_bits[317],match_bits[318],match_bits[319]});
	assign or_o[2][20]=|({match_bits[324],match_bits[325],match_bits[326],match_bits[327],match_bits[332],match_bits[333],match_bits[334],match_bits[335]});
	assign or_o[2][21]=|({match_bits[340],match_bits[341],match_bits[342],match_bits[343],match_bits[348],match_bits[349],match_bits[350],match_bits[351]});
	assign or_o[2][22]=|({match_bits[356],match_bits[357],match_bits[358],match_bits[359],match_bits[364],match_bits[365],match_bits[366],match_bits[367]});
	assign or_o[2][23]=|({match_bits[372],match_bits[373],match_bits[374],match_bits[375],match_bits[380],match_bits[381],match_bits[382],match_bits[383]});
	assign or_o[2][24]=|({match_bits[388],match_bits[389],match_bits[390],match_bits[391],match_bits[396],match_bits[397],match_bits[398],match_bits[399]});
	assign or_o[2][25]=|({match_bits[404],match_bits[405],match_bits[406],match_bits[407],match_bits[412],match_bits[413],match_bits[414],match_bits[415]});
	assign or_o[2][26]=|({match_bits[420],match_bits[421],match_bits[422],match_bits[423],match_bits[428],match_bits[429],match_bits[430],match_bits[431]});
	assign or_o[2][27]=|({match_bits[436],match_bits[437],match_bits[438],match_bits[439],match_bits[444],match_bits[445],match_bits[446],match_bits[447]});
	assign or_o[2][28]=|({match_bits[452],match_bits[453],match_bits[454],match_bits[455],match_bits[460],match_bits[461],match_bits[462],match_bits[463]});
	assign or_o[2][29]=|({match_bits[468],match_bits[469],match_bits[470],match_bits[471],match_bits[476],match_bits[477],match_bits[478],match_bits[479]});
	assign or_o[2][30]=|({match_bits[484],match_bits[485],match_bits[486],match_bits[487],match_bits[492],match_bits[493],match_bits[494],match_bits[495]});
	assign or_o[2][31]=|({match_bits[500],match_bits[501],match_bits[502],match_bits[503],match_bits[508],match_bits[509],match_bits[510],match_bits[511]});
	assign match_index[2]=|({or_o[2][0],or_o[2][1],or_o[2][2],or_o[2][3],or_o[2][4],or_o[2][5],or_o[2][6],or_o[2][7],or_o[2][8],or_o[2][9],or_o[2][10],or_o[2][11],or_o[2][12],or_o[2][13],or_o[2][14],or_o[2][15],or_o[2][16],or_o[2][17],or_o[2][18],or_o[2][19],or_o[2][20],or_o[2][21],or_o[2][22],or_o[2][23],or_o[2][24],or_o[2][25],or_o[2][26],or_o[2][27],or_o[2][28],or_o[2][29],or_o[2][30],or_o[2][31]});
	assign or_o[3][0]=|({match_bits[8],match_bits[9],match_bits[10],match_bits[11],match_bits[12],match_bits[13],match_bits[14],match_bits[15]});
	assign or_o[3][1]=|({match_bits[24],match_bits[25],match_bits[26],match_bits[27],match_bits[28],match_bits[29],match_bits[30],match_bits[31]});
	assign or_o[3][2]=|({match_bits[40],match_bits[41],match_bits[42],match_bits[43],match_bits[44],match_bits[45],match_bits[46],match_bits[47]});
	assign or_o[3][3]=|({match_bits[56],match_bits[57],match_bits[58],match_bits[59],match_bits[60],match_bits[61],match_bits[62],match_bits[63]});
	assign or_o[3][4]=|({match_bits[72],match_bits[73],match_bits[74],match_bits[75],match_bits[76],match_bits[77],match_bits[78],match_bits[79]});
	assign or_o[3][5]=|({match_bits[88],match_bits[89],match_bits[90],match_bits[91],match_bits[92],match_bits[93],match_bits[94],match_bits[95]});
	assign or_o[3][6]=|({match_bits[104],match_bits[105],match_bits[106],match_bits[107],match_bits[108],match_bits[109],match_bits[110],match_bits[111]});
	assign or_o[3][7]=|({match_bits[120],match_bits[121],match_bits[122],match_bits[123],match_bits[124],match_bits[125],match_bits[126],match_bits[127]});
	assign or_o[3][8]=|({match_bits[136],match_bits[137],match_bits[138],match_bits[139],match_bits[140],match_bits[141],match_bits[142],match_bits[143]});
	assign or_o[3][9]=|({match_bits[152],match_bits[153],match_bits[154],match_bits[155],match_bits[156],match_bits[157],match_bits[158],match_bits[159]});
	assign or_o[3][10]=|({match_bits[168],match_bits[169],match_bits[170],match_bits[171],match_bits[172],match_bits[173],match_bits[174],match_bits[175]});
	assign or_o[3][11]=|({match_bits[184],match_bits[185],match_bits[186],match_bits[187],match_bits[188],match_bits[189],match_bits[190],match_bits[191]});
	assign or_o[3][12]=|({match_bits[200],match_bits[201],match_bits[202],match_bits[203],match_bits[204],match_bits[205],match_bits[206],match_bits[207]});
	assign or_o[3][13]=|({match_bits[216],match_bits[217],match_bits[218],match_bits[219],match_bits[220],match_bits[221],match_bits[222],match_bits[223]});
	assign or_o[3][14]=|({match_bits[232],match_bits[233],match_bits[234],match_bits[235],match_bits[236],match_bits[237],match_bits[238],match_bits[239]});
	assign or_o[3][15]=|({match_bits[248],match_bits[249],match_bits[250],match_bits[251],match_bits[252],match_bits[253],match_bits[254],match_bits[255]});
	assign or_o[3][16]=|({match_bits[264],match_bits[265],match_bits[266],match_bits[267],match_bits[268],match_bits[269],match_bits[270],match_bits[271]});
	assign or_o[3][17]=|({match_bits[280],match_bits[281],match_bits[282],match_bits[283],match_bits[284],match_bits[285],match_bits[286],match_bits[287]});
	assign or_o[3][18]=|({match_bits[296],match_bits[297],match_bits[298],match_bits[299],match_bits[300],match_bits[301],match_bits[302],match_bits[303]});
	assign or_o[3][19]=|({match_bits[312],match_bits[313],match_bits[314],match_bits[315],match_bits[316],match_bits[317],match_bits[318],match_bits[319]});
	assign or_o[3][20]=|({match_bits[328],match_bits[329],match_bits[330],match_bits[331],match_bits[332],match_bits[333],match_bits[334],match_bits[335]});
	assign or_o[3][21]=|({match_bits[344],match_bits[345],match_bits[346],match_bits[347],match_bits[348],match_bits[349],match_bits[350],match_bits[351]});
	assign or_o[3][22]=|({match_bits[360],match_bits[361],match_bits[362],match_bits[363],match_bits[364],match_bits[365],match_bits[366],match_bits[367]});
	assign or_o[3][23]=|({match_bits[376],match_bits[377],match_bits[378],match_bits[379],match_bits[380],match_bits[381],match_bits[382],match_bits[383]});
	assign or_o[3][24]=|({match_bits[392],match_bits[393],match_bits[394],match_bits[395],match_bits[396],match_bits[397],match_bits[398],match_bits[399]});
	assign or_o[3][25]=|({match_bits[408],match_bits[409],match_bits[410],match_bits[411],match_bits[412],match_bits[413],match_bits[414],match_bits[415]});
	assign or_o[3][26]=|({match_bits[424],match_bits[425],match_bits[426],match_bits[427],match_bits[428],match_bits[429],match_bits[430],match_bits[431]});
	assign or_o[3][27]=|({match_bits[440],match_bits[441],match_bits[442],match_bits[443],match_bits[444],match_bits[445],match_bits[446],match_bits[447]});
	assign or_o[3][28]=|({match_bits[456],match_bits[457],match_bits[458],match_bits[459],match_bits[460],match_bits[461],match_bits[462],match_bits[463]});
	assign or_o[3][29]=|({match_bits[472],match_bits[473],match_bits[474],match_bits[475],match_bits[476],match_bits[477],match_bits[478],match_bits[479]});
	assign or_o[3][30]=|({match_bits[488],match_bits[489],match_bits[490],match_bits[491],match_bits[492],match_bits[493],match_bits[494],match_bits[495]});
	assign or_o[3][31]=|({match_bits[504],match_bits[505],match_bits[506],match_bits[507],match_bits[508],match_bits[509],match_bits[510],match_bits[511]});
	assign match_index[3]=|({or_o[3][0],or_o[3][1],or_o[3][2],or_o[3][3],or_o[3][4],or_o[3][5],or_o[3][6],or_o[3][7],or_o[3][8],or_o[3][9],or_o[3][10],or_o[3][11],or_o[3][12],or_o[3][13],or_o[3][14],or_o[3][15],or_o[3][16],or_o[3][17],or_o[3][18],or_o[3][19],or_o[3][20],or_o[3][21],or_o[3][22],or_o[3][23],or_o[3][24],or_o[3][25],or_o[3][26],or_o[3][27],or_o[3][28],or_o[3][29],or_o[3][30],or_o[3][31]});
	assign or_o[4][0]=|({match_bits[16],match_bits[17],match_bits[18],match_bits[19],match_bits[20],match_bits[21],match_bits[22],match_bits[23]});
	assign or_o[4][1]=|({match_bits[24],match_bits[25],match_bits[26],match_bits[27],match_bits[28],match_bits[29],match_bits[30],match_bits[31]});
	assign or_o[4][2]=|({match_bits[48],match_bits[49],match_bits[50],match_bits[51],match_bits[52],match_bits[53],match_bits[54],match_bits[55]});
	assign or_o[4][3]=|({match_bits[56],match_bits[57],match_bits[58],match_bits[59],match_bits[60],match_bits[61],match_bits[62],match_bits[63]});
	assign or_o[4][4]=|({match_bits[80],match_bits[81],match_bits[82],match_bits[83],match_bits[84],match_bits[85],match_bits[86],match_bits[87]});
	assign or_o[4][5]=|({match_bits[88],match_bits[89],match_bits[90],match_bits[91],match_bits[92],match_bits[93],match_bits[94],match_bits[95]});
	assign or_o[4][6]=|({match_bits[112],match_bits[113],match_bits[114],match_bits[115],match_bits[116],match_bits[117],match_bits[118],match_bits[119]});
	assign or_o[4][7]=|({match_bits[120],match_bits[121],match_bits[122],match_bits[123],match_bits[124],match_bits[125],match_bits[126],match_bits[127]});
	assign or_o[4][8]=|({match_bits[144],match_bits[145],match_bits[146],match_bits[147],match_bits[148],match_bits[149],match_bits[150],match_bits[151]});
	assign or_o[4][9]=|({match_bits[152],match_bits[153],match_bits[154],match_bits[155],match_bits[156],match_bits[157],match_bits[158],match_bits[159]});
	assign or_o[4][10]=|({match_bits[176],match_bits[177],match_bits[178],match_bits[179],match_bits[180],match_bits[181],match_bits[182],match_bits[183]});
	assign or_o[4][11]=|({match_bits[184],match_bits[185],match_bits[186],match_bits[187],match_bits[188],match_bits[189],match_bits[190],match_bits[191]});
	assign or_o[4][12]=|({match_bits[208],match_bits[209],match_bits[210],match_bits[211],match_bits[212],match_bits[213],match_bits[214],match_bits[215]});
	assign or_o[4][13]=|({match_bits[216],match_bits[217],match_bits[218],match_bits[219],match_bits[220],match_bits[221],match_bits[222],match_bits[223]});
	assign or_o[4][14]=|({match_bits[240],match_bits[241],match_bits[242],match_bits[243],match_bits[244],match_bits[245],match_bits[246],match_bits[247]});
	assign or_o[4][15]=|({match_bits[248],match_bits[249],match_bits[250],match_bits[251],match_bits[252],match_bits[253],match_bits[254],match_bits[255]});
	assign or_o[4][16]=|({match_bits[272],match_bits[273],match_bits[274],match_bits[275],match_bits[276],match_bits[277],match_bits[278],match_bits[279]});
	assign or_o[4][17]=|({match_bits[280],match_bits[281],match_bits[282],match_bits[283],match_bits[284],match_bits[285],match_bits[286],match_bits[287]});
	assign or_o[4][18]=|({match_bits[304],match_bits[305],match_bits[306],match_bits[307],match_bits[308],match_bits[309],match_bits[310],match_bits[311]});
	assign or_o[4][19]=|({match_bits[312],match_bits[313],match_bits[314],match_bits[315],match_bits[316],match_bits[317],match_bits[318],match_bits[319]});
	assign or_o[4][20]=|({match_bits[336],match_bits[337],match_bits[338],match_bits[339],match_bits[340],match_bits[341],match_bits[342],match_bits[343]});
	assign or_o[4][21]=|({match_bits[344],match_bits[345],match_bits[346],match_bits[347],match_bits[348],match_bits[349],match_bits[350],match_bits[351]});
	assign or_o[4][22]=|({match_bits[368],match_bits[369],match_bits[370],match_bits[371],match_bits[372],match_bits[373],match_bits[374],match_bits[375]});
	assign or_o[4][23]=|({match_bits[376],match_bits[377],match_bits[378],match_bits[379],match_bits[380],match_bits[381],match_bits[382],match_bits[383]});
	assign or_o[4][24]=|({match_bits[400],match_bits[401],match_bits[402],match_bits[403],match_bits[404],match_bits[405],match_bits[406],match_bits[407]});
	assign or_o[4][25]=|({match_bits[408],match_bits[409],match_bits[410],match_bits[411],match_bits[412],match_bits[413],match_bits[414],match_bits[415]});
	assign or_o[4][26]=|({match_bits[432],match_bits[433],match_bits[434],match_bits[435],match_bits[436],match_bits[437],match_bits[438],match_bits[439]});
	assign or_o[4][27]=|({match_bits[440],match_bits[441],match_bits[442],match_bits[443],match_bits[444],match_bits[445],match_bits[446],match_bits[447]});
	assign or_o[4][28]=|({match_bits[464],match_bits[465],match_bits[466],match_bits[467],match_bits[468],match_bits[469],match_bits[470],match_bits[471]});
	assign or_o[4][29]=|({match_bits[472],match_bits[473],match_bits[474],match_bits[475],match_bits[476],match_bits[477],match_bits[478],match_bits[479]});
	assign or_o[4][30]=|({match_bits[496],match_bits[497],match_bits[498],match_bits[499],match_bits[500],match_bits[501],match_bits[502],match_bits[503]});
	assign or_o[4][31]=|({match_bits[504],match_bits[505],match_bits[506],match_bits[507],match_bits[508],match_bits[509],match_bits[510],match_bits[511]});
	assign match_index[4]=|({or_o[4][0],or_o[4][1],or_o[4][2],or_o[4][3],or_o[4][4],or_o[4][5],or_o[4][6],or_o[4][7],or_o[4][8],or_o[4][9],or_o[4][10],or_o[4][11],or_o[4][12],or_o[4][13],or_o[4][14],or_o[4][15],or_o[4][16],or_o[4][17],or_o[4][18],or_o[4][19],or_o[4][20],or_o[4][21],or_o[4][22],or_o[4][23],or_o[4][24],or_o[4][25],or_o[4][26],or_o[4][27],or_o[4][28],or_o[4][29],or_o[4][30],or_o[4][31]});
	assign or_o[5][0]=|({match_bits[32],match_bits[33],match_bits[34],match_bits[35],match_bits[36],match_bits[37],match_bits[38],match_bits[39]});
	assign or_o[5][1]=|({match_bits[40],match_bits[41],match_bits[42],match_bits[43],match_bits[44],match_bits[45],match_bits[46],match_bits[47]});
	assign or_o[5][2]=|({match_bits[48],match_bits[49],match_bits[50],match_bits[51],match_bits[52],match_bits[53],match_bits[54],match_bits[55]});
	assign or_o[5][3]=|({match_bits[56],match_bits[57],match_bits[58],match_bits[59],match_bits[60],match_bits[61],match_bits[62],match_bits[63]});
	assign or_o[5][4]=|({match_bits[96],match_bits[97],match_bits[98],match_bits[99],match_bits[100],match_bits[101],match_bits[102],match_bits[103]});
	assign or_o[5][5]=|({match_bits[104],match_bits[105],match_bits[106],match_bits[107],match_bits[108],match_bits[109],match_bits[110],match_bits[111]});
	assign or_o[5][6]=|({match_bits[112],match_bits[113],match_bits[114],match_bits[115],match_bits[116],match_bits[117],match_bits[118],match_bits[119]});
	assign or_o[5][7]=|({match_bits[120],match_bits[121],match_bits[122],match_bits[123],match_bits[124],match_bits[125],match_bits[126],match_bits[127]});
	assign or_o[5][8]=|({match_bits[160],match_bits[161],match_bits[162],match_bits[163],match_bits[164],match_bits[165],match_bits[166],match_bits[167]});
	assign or_o[5][9]=|({match_bits[168],match_bits[169],match_bits[170],match_bits[171],match_bits[172],match_bits[173],match_bits[174],match_bits[175]});
	assign or_o[5][10]=|({match_bits[176],match_bits[177],match_bits[178],match_bits[179],match_bits[180],match_bits[181],match_bits[182],match_bits[183]});
	assign or_o[5][11]=|({match_bits[184],match_bits[185],match_bits[186],match_bits[187],match_bits[188],match_bits[189],match_bits[190],match_bits[191]});
	assign or_o[5][12]=|({match_bits[224],match_bits[225],match_bits[226],match_bits[227],match_bits[228],match_bits[229],match_bits[230],match_bits[231]});
	assign or_o[5][13]=|({match_bits[232],match_bits[233],match_bits[234],match_bits[235],match_bits[236],match_bits[237],match_bits[238],match_bits[239]});
	assign or_o[5][14]=|({match_bits[240],match_bits[241],match_bits[242],match_bits[243],match_bits[244],match_bits[245],match_bits[246],match_bits[247]});
	assign or_o[5][15]=|({match_bits[248],match_bits[249],match_bits[250],match_bits[251],match_bits[252],match_bits[253],match_bits[254],match_bits[255]});
	assign or_o[5][16]=|({match_bits[288],match_bits[289],match_bits[290],match_bits[291],match_bits[292],match_bits[293],match_bits[294],match_bits[295]});
	assign or_o[5][17]=|({match_bits[296],match_bits[297],match_bits[298],match_bits[299],match_bits[300],match_bits[301],match_bits[302],match_bits[303]});
	assign or_o[5][18]=|({match_bits[304],match_bits[305],match_bits[306],match_bits[307],match_bits[308],match_bits[309],match_bits[310],match_bits[311]});
	assign or_o[5][19]=|({match_bits[312],match_bits[313],match_bits[314],match_bits[315],match_bits[316],match_bits[317],match_bits[318],match_bits[319]});
	assign or_o[5][20]=|({match_bits[352],match_bits[353],match_bits[354],match_bits[355],match_bits[356],match_bits[357],match_bits[358],match_bits[359]});
	assign or_o[5][21]=|({match_bits[360],match_bits[361],match_bits[362],match_bits[363],match_bits[364],match_bits[365],match_bits[366],match_bits[367]});
	assign or_o[5][22]=|({match_bits[368],match_bits[369],match_bits[370],match_bits[371],match_bits[372],match_bits[373],match_bits[374],match_bits[375]});
	assign or_o[5][23]=|({match_bits[376],match_bits[377],match_bits[378],match_bits[379],match_bits[380],match_bits[381],match_bits[382],match_bits[383]});
	assign or_o[5][24]=|({match_bits[416],match_bits[417],match_bits[418],match_bits[419],match_bits[420],match_bits[421],match_bits[422],match_bits[423]});
	assign or_o[5][25]=|({match_bits[424],match_bits[425],match_bits[426],match_bits[427],match_bits[428],match_bits[429],match_bits[430],match_bits[431]});
	assign or_o[5][26]=|({match_bits[432],match_bits[433],match_bits[434],match_bits[435],match_bits[436],match_bits[437],match_bits[438],match_bits[439]});
	assign or_o[5][27]=|({match_bits[440],match_bits[441],match_bits[442],match_bits[443],match_bits[444],match_bits[445],match_bits[446],match_bits[447]});
	assign or_o[5][28]=|({match_bits[480],match_bits[481],match_bits[482],match_bits[483],match_bits[484],match_bits[485],match_bits[486],match_bits[487]});
	assign or_o[5][29]=|({match_bits[488],match_bits[489],match_bits[490],match_bits[491],match_bits[492],match_bits[493],match_bits[494],match_bits[495]});
	assign or_o[5][30]=|({match_bits[496],match_bits[497],match_bits[498],match_bits[499],match_bits[500],match_bits[501],match_bits[502],match_bits[503]});
	assign or_o[5][31]=|({match_bits[504],match_bits[505],match_bits[506],match_bits[507],match_bits[508],match_bits[509],match_bits[510],match_bits[511]});
	assign match_index[5]=|({or_o[5][0],or_o[5][1],or_o[5][2],or_o[5][3],or_o[5][4],or_o[5][5],or_o[5][6],or_o[5][7],or_o[5][8],or_o[5][9],or_o[5][10],or_o[5][11],or_o[5][12],or_o[5][13],or_o[5][14],or_o[5][15],or_o[5][16],or_o[5][17],or_o[5][18],or_o[5][19],or_o[5][20],or_o[5][21],or_o[5][22],or_o[5][23],or_o[5][24],or_o[5][25],or_o[5][26],or_o[5][27],or_o[5][28],or_o[5][29],or_o[5][30],or_o[5][31]});
	assign or_o[6][0]=|({match_bits[64],match_bits[65],match_bits[66],match_bits[67],match_bits[68],match_bits[69],match_bits[70],match_bits[71]});
	assign or_o[6][1]=|({match_bits[72],match_bits[73],match_bits[74],match_bits[75],match_bits[76],match_bits[77],match_bits[78],match_bits[79]});
	assign or_o[6][2]=|({match_bits[80],match_bits[81],match_bits[82],match_bits[83],match_bits[84],match_bits[85],match_bits[86],match_bits[87]});
	assign or_o[6][3]=|({match_bits[88],match_bits[89],match_bits[90],match_bits[91],match_bits[92],match_bits[93],match_bits[94],match_bits[95]});
	assign or_o[6][4]=|({match_bits[96],match_bits[97],match_bits[98],match_bits[99],match_bits[100],match_bits[101],match_bits[102],match_bits[103]});
	assign or_o[6][5]=|({match_bits[104],match_bits[105],match_bits[106],match_bits[107],match_bits[108],match_bits[109],match_bits[110],match_bits[111]});
	assign or_o[6][6]=|({match_bits[112],match_bits[113],match_bits[114],match_bits[115],match_bits[116],match_bits[117],match_bits[118],match_bits[119]});
	assign or_o[6][7]=|({match_bits[120],match_bits[121],match_bits[122],match_bits[123],match_bits[124],match_bits[125],match_bits[126],match_bits[127]});
	assign or_o[6][8]=|({match_bits[192],match_bits[193],match_bits[194],match_bits[195],match_bits[196],match_bits[197],match_bits[198],match_bits[199]});
	assign or_o[6][9]=|({match_bits[200],match_bits[201],match_bits[202],match_bits[203],match_bits[204],match_bits[205],match_bits[206],match_bits[207]});
	assign or_o[6][10]=|({match_bits[208],match_bits[209],match_bits[210],match_bits[211],match_bits[212],match_bits[213],match_bits[214],match_bits[215]});
	assign or_o[6][11]=|({match_bits[216],match_bits[217],match_bits[218],match_bits[219],match_bits[220],match_bits[221],match_bits[222],match_bits[223]});
	assign or_o[6][12]=|({match_bits[224],match_bits[225],match_bits[226],match_bits[227],match_bits[228],match_bits[229],match_bits[230],match_bits[231]});
	assign or_o[6][13]=|({match_bits[232],match_bits[233],match_bits[234],match_bits[235],match_bits[236],match_bits[237],match_bits[238],match_bits[239]});
	assign or_o[6][14]=|({match_bits[240],match_bits[241],match_bits[242],match_bits[243],match_bits[244],match_bits[245],match_bits[246],match_bits[247]});
	assign or_o[6][15]=|({match_bits[248],match_bits[249],match_bits[250],match_bits[251],match_bits[252],match_bits[253],match_bits[254],match_bits[255]});
	assign or_o[6][16]=|({match_bits[320],match_bits[321],match_bits[322],match_bits[323],match_bits[324],match_bits[325],match_bits[326],match_bits[327]});
	assign or_o[6][17]=|({match_bits[328],match_bits[329],match_bits[330],match_bits[331],match_bits[332],match_bits[333],match_bits[334],match_bits[335]});
	assign or_o[6][18]=|({match_bits[336],match_bits[337],match_bits[338],match_bits[339],match_bits[340],match_bits[341],match_bits[342],match_bits[343]});
	assign or_o[6][19]=|({match_bits[344],match_bits[345],match_bits[346],match_bits[347],match_bits[348],match_bits[349],match_bits[350],match_bits[351]});
	assign or_o[6][20]=|({match_bits[352],match_bits[353],match_bits[354],match_bits[355],match_bits[356],match_bits[357],match_bits[358],match_bits[359]});
	assign or_o[6][21]=|({match_bits[360],match_bits[361],match_bits[362],match_bits[363],match_bits[364],match_bits[365],match_bits[366],match_bits[367]});
	assign or_o[6][22]=|({match_bits[368],match_bits[369],match_bits[370],match_bits[371],match_bits[372],match_bits[373],match_bits[374],match_bits[375]});
	assign or_o[6][23]=|({match_bits[376],match_bits[377],match_bits[378],match_bits[379],match_bits[380],match_bits[381],match_bits[382],match_bits[383]});
	assign or_o[6][24]=|({match_bits[448],match_bits[449],match_bits[450],match_bits[451],match_bits[452],match_bits[453],match_bits[454],match_bits[455]});
	assign or_o[6][25]=|({match_bits[456],match_bits[457],match_bits[458],match_bits[459],match_bits[460],match_bits[461],match_bits[462],match_bits[463]});
	assign or_o[6][26]=|({match_bits[464],match_bits[465],match_bits[466],match_bits[467],match_bits[468],match_bits[469],match_bits[470],match_bits[471]});
	assign or_o[6][27]=|({match_bits[472],match_bits[473],match_bits[474],match_bits[475],match_bits[476],match_bits[477],match_bits[478],match_bits[479]});
	assign or_o[6][28]=|({match_bits[480],match_bits[481],match_bits[482],match_bits[483],match_bits[484],match_bits[485],match_bits[486],match_bits[487]});
	assign or_o[6][29]=|({match_bits[488],match_bits[489],match_bits[490],match_bits[491],match_bits[492],match_bits[493],match_bits[494],match_bits[495]});
	assign or_o[6][30]=|({match_bits[496],match_bits[497],match_bits[498],match_bits[499],match_bits[500],match_bits[501],match_bits[502],match_bits[503]});
	assign or_o[6][31]=|({match_bits[504],match_bits[505],match_bits[506],match_bits[507],match_bits[508],match_bits[509],match_bits[510],match_bits[511]});
	assign match_index[6]=|({or_o[6][0],or_o[6][1],or_o[6][2],or_o[6][3],or_o[6][4],or_o[6][5],or_o[6][6],or_o[6][7],or_o[6][8],or_o[6][9],or_o[6][10],or_o[6][11],or_o[6][12],or_o[6][13],or_o[6][14],or_o[6][15],or_o[6][16],or_o[6][17],or_o[6][18],or_o[6][19],or_o[6][20],or_o[6][21],or_o[6][22],or_o[6][23],or_o[6][24],or_o[6][25],or_o[6][26],or_o[6][27],or_o[6][28],or_o[6][29],or_o[6][30],or_o[6][31]});
	assign or_o[7][0]=|({match_bits[128],match_bits[129],match_bits[130],match_bits[131],match_bits[132],match_bits[133],match_bits[134],match_bits[135]});
	assign or_o[7][1]=|({match_bits[136],match_bits[137],match_bits[138],match_bits[139],match_bits[140],match_bits[141],match_bits[142],match_bits[143]});
	assign or_o[7][2]=|({match_bits[144],match_bits[145],match_bits[146],match_bits[147],match_bits[148],match_bits[149],match_bits[150],match_bits[151]});
	assign or_o[7][3]=|({match_bits[152],match_bits[153],match_bits[154],match_bits[155],match_bits[156],match_bits[157],match_bits[158],match_bits[159]});
	assign or_o[7][4]=|({match_bits[160],match_bits[161],match_bits[162],match_bits[163],match_bits[164],match_bits[165],match_bits[166],match_bits[167]});
	assign or_o[7][5]=|({match_bits[168],match_bits[169],match_bits[170],match_bits[171],match_bits[172],match_bits[173],match_bits[174],match_bits[175]});
	assign or_o[7][6]=|({match_bits[176],match_bits[177],match_bits[178],match_bits[179],match_bits[180],match_bits[181],match_bits[182],match_bits[183]});
	assign or_o[7][7]=|({match_bits[184],match_bits[185],match_bits[186],match_bits[187],match_bits[188],match_bits[189],match_bits[190],match_bits[191]});
	assign or_o[7][8]=|({match_bits[192],match_bits[193],match_bits[194],match_bits[195],match_bits[196],match_bits[197],match_bits[198],match_bits[199]});
	assign or_o[7][9]=|({match_bits[200],match_bits[201],match_bits[202],match_bits[203],match_bits[204],match_bits[205],match_bits[206],match_bits[207]});
	assign or_o[7][10]=|({match_bits[208],match_bits[209],match_bits[210],match_bits[211],match_bits[212],match_bits[213],match_bits[214],match_bits[215]});
	assign or_o[7][11]=|({match_bits[216],match_bits[217],match_bits[218],match_bits[219],match_bits[220],match_bits[221],match_bits[222],match_bits[223]});
	assign or_o[7][12]=|({match_bits[224],match_bits[225],match_bits[226],match_bits[227],match_bits[228],match_bits[229],match_bits[230],match_bits[231]});
	assign or_o[7][13]=|({match_bits[232],match_bits[233],match_bits[234],match_bits[235],match_bits[236],match_bits[237],match_bits[238],match_bits[239]});
	assign or_o[7][14]=|({match_bits[240],match_bits[241],match_bits[242],match_bits[243],match_bits[244],match_bits[245],match_bits[246],match_bits[247]});
	assign or_o[7][15]=|({match_bits[248],match_bits[249],match_bits[250],match_bits[251],match_bits[252],match_bits[253],match_bits[254],match_bits[255]});
	assign or_o[7][16]=|({match_bits[384],match_bits[385],match_bits[386],match_bits[387],match_bits[388],match_bits[389],match_bits[390],match_bits[391]});
	assign or_o[7][17]=|({match_bits[392],match_bits[393],match_bits[394],match_bits[395],match_bits[396],match_bits[397],match_bits[398],match_bits[399]});
	assign or_o[7][18]=|({match_bits[400],match_bits[401],match_bits[402],match_bits[403],match_bits[404],match_bits[405],match_bits[406],match_bits[407]});
	assign or_o[7][19]=|({match_bits[408],match_bits[409],match_bits[410],match_bits[411],match_bits[412],match_bits[413],match_bits[414],match_bits[415]});
	assign or_o[7][20]=|({match_bits[416],match_bits[417],match_bits[418],match_bits[419],match_bits[420],match_bits[421],match_bits[422],match_bits[423]});
	assign or_o[7][21]=|({match_bits[424],match_bits[425],match_bits[426],match_bits[427],match_bits[428],match_bits[429],match_bits[430],match_bits[431]});
	assign or_o[7][22]=|({match_bits[432],match_bits[433],match_bits[434],match_bits[435],match_bits[436],match_bits[437],match_bits[438],match_bits[439]});
	assign or_o[7][23]=|({match_bits[440],match_bits[441],match_bits[442],match_bits[443],match_bits[444],match_bits[445],match_bits[446],match_bits[447]});
	assign or_o[7][24]=|({match_bits[448],match_bits[449],match_bits[450],match_bits[451],match_bits[452],match_bits[453],match_bits[454],match_bits[455]});
	assign or_o[7][25]=|({match_bits[456],match_bits[457],match_bits[458],match_bits[459],match_bits[460],match_bits[461],match_bits[462],match_bits[463]});
	assign or_o[7][26]=|({match_bits[464],match_bits[465],match_bits[466],match_bits[467],match_bits[468],match_bits[469],match_bits[470],match_bits[471]});
	assign or_o[7][27]=|({match_bits[472],match_bits[473],match_bits[474],match_bits[475],match_bits[476],match_bits[477],match_bits[478],match_bits[479]});
	assign or_o[7][28]=|({match_bits[480],match_bits[481],match_bits[482],match_bits[483],match_bits[484],match_bits[485],match_bits[486],match_bits[487]});
	assign or_o[7][29]=|({match_bits[488],match_bits[489],match_bits[490],match_bits[491],match_bits[492],match_bits[493],match_bits[494],match_bits[495]});
	assign or_o[7][30]=|({match_bits[496],match_bits[497],match_bits[498],match_bits[499],match_bits[500],match_bits[501],match_bits[502],match_bits[503]});
	assign or_o[7][31]=|({match_bits[504],match_bits[505],match_bits[506],match_bits[507],match_bits[508],match_bits[509],match_bits[510],match_bits[511]});
	assign match_index[7]=|({or_o[7][0],or_o[7][1],or_o[7][2],or_o[7][3],or_o[7][4],or_o[7][5],or_o[7][6],or_o[7][7],or_o[7][8],or_o[7][9],or_o[7][10],or_o[7][11],or_o[7][12],or_o[7][13],or_o[7][14],or_o[7][15],or_o[7][16],or_o[7][17],or_o[7][18],or_o[7][19],or_o[7][20],or_o[7][21],or_o[7][22],or_o[7][23],or_o[7][24],or_o[7][25],or_o[7][26],or_o[7][27],or_o[7][28],or_o[7][29],or_o[7][30],or_o[7][31]});
	assign or_o[8][0]=|({match_bits[256],match_bits[257],match_bits[258],match_bits[259],match_bits[260],match_bits[261],match_bits[262],match_bits[263]});
	assign or_o[8][1]=|({match_bits[264],match_bits[265],match_bits[266],match_bits[267],match_bits[268],match_bits[269],match_bits[270],match_bits[271]});
	assign or_o[8][2]=|({match_bits[272],match_bits[273],match_bits[274],match_bits[275],match_bits[276],match_bits[277],match_bits[278],match_bits[279]});
	assign or_o[8][3]=|({match_bits[280],match_bits[281],match_bits[282],match_bits[283],match_bits[284],match_bits[285],match_bits[286],match_bits[287]});
	assign or_o[8][4]=|({match_bits[288],match_bits[289],match_bits[290],match_bits[291],match_bits[292],match_bits[293],match_bits[294],match_bits[295]});
	assign or_o[8][5]=|({match_bits[296],match_bits[297],match_bits[298],match_bits[299],match_bits[300],match_bits[301],match_bits[302],match_bits[303]});
	assign or_o[8][6]=|({match_bits[304],match_bits[305],match_bits[306],match_bits[307],match_bits[308],match_bits[309],match_bits[310],match_bits[311]});
	assign or_o[8][7]=|({match_bits[312],match_bits[313],match_bits[314],match_bits[315],match_bits[316],match_bits[317],match_bits[318],match_bits[319]});
	assign or_o[8][8]=|({match_bits[320],match_bits[321],match_bits[322],match_bits[323],match_bits[324],match_bits[325],match_bits[326],match_bits[327]});
	assign or_o[8][9]=|({match_bits[328],match_bits[329],match_bits[330],match_bits[331],match_bits[332],match_bits[333],match_bits[334],match_bits[335]});
	assign or_o[8][10]=|({match_bits[336],match_bits[337],match_bits[338],match_bits[339],match_bits[340],match_bits[341],match_bits[342],match_bits[343]});
	assign or_o[8][11]=|({match_bits[344],match_bits[345],match_bits[346],match_bits[347],match_bits[348],match_bits[349],match_bits[350],match_bits[351]});
	assign or_o[8][12]=|({match_bits[352],match_bits[353],match_bits[354],match_bits[355],match_bits[356],match_bits[357],match_bits[358],match_bits[359]});
	assign or_o[8][13]=|({match_bits[360],match_bits[361],match_bits[362],match_bits[363],match_bits[364],match_bits[365],match_bits[366],match_bits[367]});
	assign or_o[8][14]=|({match_bits[368],match_bits[369],match_bits[370],match_bits[371],match_bits[372],match_bits[373],match_bits[374],match_bits[375]});
	assign or_o[8][15]=|({match_bits[376],match_bits[377],match_bits[378],match_bits[379],match_bits[380],match_bits[381],match_bits[382],match_bits[383]});
	assign or_o[8][16]=|({match_bits[384],match_bits[385],match_bits[386],match_bits[387],match_bits[388],match_bits[389],match_bits[390],match_bits[391]});
	assign or_o[8][17]=|({match_bits[392],match_bits[393],match_bits[394],match_bits[395],match_bits[396],match_bits[397],match_bits[398],match_bits[399]});
	assign or_o[8][18]=|({match_bits[400],match_bits[401],match_bits[402],match_bits[403],match_bits[404],match_bits[405],match_bits[406],match_bits[407]});
	assign or_o[8][19]=|({match_bits[408],match_bits[409],match_bits[410],match_bits[411],match_bits[412],match_bits[413],match_bits[414],match_bits[415]});
	assign or_o[8][20]=|({match_bits[416],match_bits[417],match_bits[418],match_bits[419],match_bits[420],match_bits[421],match_bits[422],match_bits[423]});
	assign or_o[8][21]=|({match_bits[424],match_bits[425],match_bits[426],match_bits[427],match_bits[428],match_bits[429],match_bits[430],match_bits[431]});
	assign or_o[8][22]=|({match_bits[432],match_bits[433],match_bits[434],match_bits[435],match_bits[436],match_bits[437],match_bits[438],match_bits[439]});
	assign or_o[8][23]=|({match_bits[440],match_bits[441],match_bits[442],match_bits[443],match_bits[444],match_bits[445],match_bits[446],match_bits[447]});
	assign or_o[8][24]=|({match_bits[448],match_bits[449],match_bits[450],match_bits[451],match_bits[452],match_bits[453],match_bits[454],match_bits[455]});
	assign or_o[8][25]=|({match_bits[456],match_bits[457],match_bits[458],match_bits[459],match_bits[460],match_bits[461],match_bits[462],match_bits[463]});
	assign or_o[8][26]=|({match_bits[464],match_bits[465],match_bits[466],match_bits[467],match_bits[468],match_bits[469],match_bits[470],match_bits[471]});
	assign or_o[8][27]=|({match_bits[472],match_bits[473],match_bits[474],match_bits[475],match_bits[476],match_bits[477],match_bits[478],match_bits[479]});
	assign or_o[8][28]=|({match_bits[480],match_bits[481],match_bits[482],match_bits[483],match_bits[484],match_bits[485],match_bits[486],match_bits[487]});
	assign or_o[8][29]=|({match_bits[488],match_bits[489],match_bits[490],match_bits[491],match_bits[492],match_bits[493],match_bits[494],match_bits[495]});
	assign or_o[8][30]=|({match_bits[496],match_bits[497],match_bits[498],match_bits[499],match_bits[500],match_bits[501],match_bits[502],match_bits[503]});
	assign or_o[8][31]=|({match_bits[504],match_bits[505],match_bits[506],match_bits[507],match_bits[508],match_bits[509],match_bits[510],match_bits[511]});
	assign match_index[8]=|({or_o[8][0],or_o[8][1],or_o[8][2],or_o[8][3],or_o[8][4],or_o[8][5],or_o[8][6],or_o[8][7],or_o[8][8],or_o[8][9],or_o[8][10],or_o[8][11],or_o[8][12],or_o[8][13],or_o[8][14],or_o[8][15],or_o[8][16],or_o[8][17],or_o[8][18],or_o[8][19],or_o[8][20],or_o[8][21],or_o[8][22],or_o[8][23],or_o[8][24],or_o[8][25],or_o[8][26],or_o[8][27],or_o[8][28],or_o[8][29],or_o[8][30],or_o[8][31]});
always@(match_index)begin
	match_index_reg=match_index;
	actual_match=|({match_index,match_bits[0]});
end

endmodule